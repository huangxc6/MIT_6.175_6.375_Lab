// Return Address Stack

