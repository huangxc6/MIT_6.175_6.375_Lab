import Types::*;
import ProcTypes::*;
import RegFile::*;
import Vector::*;

// indexSize is the number of bits in the index
// tagSize is the number of bits in the tag
interface Btb#(numeric type indexSize, numeric type tagSize);
    method Addr predPc(Addr pc);
    method Action update(Addr thispc, Addr nextpc);
endinterface

// BTB
module mkBtb( Btb#(indexSize, tagSize) ) provisos (Add#(indexSize,a__,32), Add#(tagSize,b__,32), Add#(TAdd#(indexSize,tagSize),c__,30));
    Vector#(TExp#(indexSize), Reg#(Addr))          targets <- replicateM(mkReg(0));
    Vector#(TExp#(indexSize), Reg#(Bit#(tagSize)))    tags <- replicateM(mkReg(0));
    Vector#(TExp#(indexSize), Reg#(Bool))            valid <- replicateM(mkReg(False));

    function Bit#(indexSize) getIndex(Addr pc) = truncate(pc >> 2);
    function Bit#(tagSize) getTag(Addr pc) = truncate(pc >> (2 + valueOf(indexSize)));

    method Addr predPc(Addr pc);
        let index = getIndex(pc);
        let tag = getTag(pc);

        if(valid[index] && (tag == tags[index])) begin
            return targets[index];
        end else begin
            return (pc + 4);
        end
    endmethod

    method Action update(Addr thisPc, Addr nextPc);
        if( nextPc != thisPc + 4 ) begin
            let index = getIndex(thisPc);
            let tag = getTag(thisPc);
            // update entry
            valid[index] <= True;
            tags[index] <= tag;
            targets[index] <= nextPc;
        end
    endmethod
endmodule

